(* EVM Contract Behavior Formalization *)
(* for Coq 8.5pl2 *)

(* Yoichi Hirai i@yoichihirai.com
   Creative Commons Attribution-ShareAlike 4.0 International License *)

(* This is just a sketch of an idea put together on a weekend.
   In the interactive theorem prover Coq, I (re)started reasoning
   about a contract’s behaviour where it can be called, returned
   from a call, and of course re-entered.

   My first example is a contract that always returns, for which I
   - wrote a specification [always_return]
   - wrote some EVM code [example1_program]
   - proved that the code satisfies the specification. [example1_spec_impl_match]

   Don’t take it seriously: I haven’t checked anything against the real implementation.

   - explore other strategies modelling the infinite process
     (an Ethereum contract goes through unlimited number of events),
   - translate more parts of the yellow paper: more instructions, and the gas economics
   - check the translation against real blockchain data
   - verify gradually more complex contracts
   - develop proof methodology.
*)

(* Gas is not considered among many things.  A contract in reality dies more often than described here. *)


(***
 *** Some basic <del>definitions</del> assumptions
 ***)

(* Here I'm being lazy and assuming that these things exist.
 * I hope these don't enable us to prove 0 = 1.
 *)


(* This module can be instantiated into some concrete ways and some more abstract ways. *)
(* A word can be a tuple of 256 booleans. *)
(* Alternatively a word can be thought of as some abstract values.
 * This would be interesting in bytecode analysis tools.
 *)
(* Many aspects of the EVM semantics do not care how words are represented. *)

Require Import NArith.
Require FMapList.
Require Import OrderedType.

Require Import Word.
Require Import ContractSem.

Require Import Cyclic.Abstract.CyclicAxioms.
Require Import Coq.Lists.List.

  Require Import ZArith.

  Require BinNums.
  Require Cyclic.ZModulo.ZModulo.

(* A useful lemma to be proven *)
Lemma addsub :
  forall x y z,
    ZModulo.add (ZModulo.sub x y) z =
    ZModulo.sub (ZModulo.add x z) y.
Proof.
  unfold ZModulo.add.
  unfold ZModulo.sub.
  intros ? ? ?.
  omega.
Qed.


Lemma addK :
  forall a b, ZModulo.sub (ZModulo.add a b) b = a.
Proof.
  unfold ZModulo.add.
  unfold ZModulo.sub.
  intros ? ?; omega.
Qed.

Lemma addC (* This lemma should not enter Word. *) :
  forall a b, ZModulo.add a b = ZModulo.add b a.
Proof.
  unfold ZModulo.add.
  intros ? ?; omega.
Qed.

Module ConcreteWord <: Word.

  Module WLEN <: Cyclic.ZModulo.ZModulo.PositiveNotOne.
    Import BinNums.

    Definition p : positive := xO (xO (xO (xO (xO (xO (xO (xO xH))))))).
    Lemma not_one : p <> 1%positive.
      unfold p.
      congruence.
    Qed.
  End WLEN.

  Module BLEN <: Cyclic.ZModulo.ZModulo.PositiveNotOne.
    Import BinNums.

    Definition p : positive := xO (xO (xO xH)).
    Lemma not_one : p <> 1%positive.
      unfold p.
      congruence.
    Qed.
  End BLEN.

  Module ALEN <: Cyclic.ZModulo.ZModulo.PositiveNotOne.
    Import BinNums.

    Definition p : positive := 160.
    Lemma not_one : p <> 1%positive.
      unfold p.
      congruence.
    Qed.
  End ALEN.

  Module W := Cyclic.ZModulo.ZModulo.ZModuloCyclicType WLEN.

  Module B := Cyclic.ZModulo.ZModulo.ZModuloCyclicType BLEN.

  Module A := Cyclic.ZModulo.ZModulo.ZModuloCyclicType ALEN.

  Definition word := W.t.

  Definition word_eq (a : W.t) (b : W.t) :=
    match ZnZ.compare a b with Eq => true | _ => false end.

  Definition word_add (a b : W.t) :=
    ZnZ.add a b.

  Arguments word_add a b /.

  Definition word_mul (a b : W.t) := ZnZ.mul a b.

  Definition word_sub := ZnZ.sub.

  Definition word_one := ZnZ.one.

  Definition word_zero := ZnZ.zero.

  Definition word_iszero := ZnZ.eq0.

  Definition word_mod := ZnZ.modulo.


  Definition word_smaller a b :=
    match ZnZ.compare a b with Lt => true | _ => false end.

  Definition word_smaller_or_eq a b :=
    match ZnZ.compare a b with Lt => true | Eq => true | Gt => false end.

  Definition word_of_N := Z.of_N.

  Definition N_of_word w := Z.to_N (ZnZ.to_Z w).

  Open Scope N_scope.
  Lemma N_of_word_of_N :
    forall (n : N), n < 10000 -> N_of_word (word_of_N n) = n.
  Proof.
    intros n nsmall.
    unfold N_of_word.
    unfold word_of_N.
    unfold ZnZ.to_Z.
    simpl.
    unfold ZModulo.to_Z.
    unfold ZModulo.wB.
    unfold WLEN.p.
    unfold DoubleType.base.
    rewrite Z.mod_small.
    { rewrite N2Z.id.
      reflexivity. }
    split.
    {
      apply N2Z.is_nonneg.
    }
    {
      eapply Z.lt_trans.
      { apply N2Z.inj_lt.
        eassumption. }
      vm_compute; auto.
    }
  Qed.

  Module WordOrdered <: OrderedType.
  (* Before using FSetList as storage,
     I need word as OrderedType *)


      Definition t := W.t.
      Definition eq a b := is_true (word_eq a b).
      Arguments eq /.

      Definition lt a b := is_true (word_smaller a b).
      Arguments lt /.


      Lemma eq_refl : forall x : t, eq x x.
      Proof.
        intro.
        unfold eq.
        unfold word_eq.
        simpl.
        rewrite ZModulo.spec_compare.
        rewrite Z.compare_refl.
        auto.
      Qed.

      Lemma eq_sym : forall x y : t, eq x y -> eq y x.
      Proof.
        intros ? ?.
        simpl.
        unfold word_eq. simpl.
        rewrite !ZModulo.spec_compare.
        rewrite <-Zcompare_antisym.
        simpl.
        set (r := (ZModulo.to_Z ALEN.p y ?= ZModulo.to_Z ALEN.p x)%Z).
        case r; unfold CompOpp; auto.
      Qed.

      Lemma eq_trans : forall x y z : t, eq x y -> eq y z -> eq x z.
      Proof.
        intros ? ? ?.
        unfold eq.
        unfold word_eq.
        simpl.
        rewrite !ZModulo.spec_compare.
        set (xy := (ZModulo.to_Z ALEN.p x ?= ZModulo.to_Z ALEN.p y)%Z).
        case_eq xy; auto; try congruence.
        unfold xy.
        rewrite Z.compare_eq_iff.
        intro H.
        rewrite H.
        auto.
      Qed.

      Lemma lt_trans : forall x y z : t, lt x y -> lt y z -> lt x z.
      Proof.
        intros x y z.
        unfold lt.
        unfold word_smaller.
        simpl.
        rewrite !ZModulo.spec_compare.
        case_eq (ZModulo.to_Z ALEN.p x ?= ZModulo.to_Z ALEN.p y)%Z; try congruence.
        case_eq (ZModulo.to_Z ALEN.p y ?= ZModulo.to_Z ALEN.p z)%Z; try congruence.
        intros H I _ _.
        erewrite (Zcompare_Lt_trans); auto; eassumption.
      Qed.

      Lemma lt_not_eq : forall x y : t, lt x y -> ~ eq x y.
      Proof.
        unfold t.
        intros x y.
        unfold lt; unfold eq.
        unfold word_smaller; unfold word_eq.
        simpl.
        case_eq (ZModulo.compare ALEN.p x y); congruence.
      Qed.

      Definition compare : forall x y : t, Compare lt eq x y.
      Proof.
        intros x y.
        unfold lt.
        case_eq (word_smaller x y); intro L.
        { apply LT; auto. }
        unfold eq.
        case_eq (word_eq x y); intro E.
        { apply EQ; auto. }
        apply GT.
        unfold word_smaller.
        unfold word_smaller in L.
        unfold word_eq in E.
        simpl in *.

        rewrite ZModulo.spec_compare in *.

        case_eq (ZModulo.to_Z ALEN.p y ?= ZModulo.to_Z ALEN.p x)%Z; try congruence.

        {
          rewrite Z.compare_eq_iff.
          intro H.
          rewrite H in E.
          rewrite Z.compare_refl in E.
          congruence.
        }
        {
          rewrite Zcompare_Gt_Lt_antisym.
          intro H.
          rewrite H in L.
          congruence.
        }
      Defined.

      Definition eq_dec : forall x y : t, {eq x y} + {~ eq x y}.
      Proof.
        unfold eq.
        intros x y.
        case (word_eq x y); [left | right]; congruence.
      Defined.

  End WordOrdered.


  Definition raw_byte := B.t.
  Inductive byte' :=
  | ByteRaw : raw_byte -> byte'
  | ByteOfWord : word -> nat -> byte'
  .
  Definition byte := byte'.

  Definition address := A.t.

  Definition address_of_word (w : word) : address := w.

  Definition address_eq a b :=
    match ZnZ.compare a b with Eq => true | _ => false end.

  Lemma address_eq_refl :
    forall a, address_eq a a = true.
  Proof.
    intro a.
    unfold address_eq.
    rewrite ZnZ.spec_compare.
    rewrite Z.compare_refl.
    reflexivity.
  Qed.

  Definition word_nth_byte (w : word) (n : nat) : byte :=
    ByteOfWord w n.

  Axiom word_of_bytes : list byte -> word.

  Open Scope list_scope.

  Import ListNotations.
  Lemma words_of_nth_bytes :
    forall w b0 b1 b2 b3 b4 b5 b6 b7 b8 b9 b10 b11 b12 b13 b14 b15 b16 b17 b18 b19 b20 b21 b22 b23 b24 b25 b26 b27 b28 b29 b30 b31,
    b0 = word_nth_byte w 0 ->
    b1 = word_nth_byte w 1 ->
    b2 = word_nth_byte w 2 ->
    b3 = word_nth_byte w 3 ->
    b4 = word_nth_byte w 4 ->
    b5 = word_nth_byte w 5 ->
    b6 = word_nth_byte w 6 ->
    b7 = word_nth_byte w 7 ->
    b8 = word_nth_byte w 8 ->
    b9 = word_nth_byte w 9 ->
    b10 = word_nth_byte w 10 ->
    b11 = word_nth_byte w 11 ->
    b12 = word_nth_byte w 12 ->
    b13 = word_nth_byte w 13 ->
    b14 = word_nth_byte w 14 ->
    b15 = word_nth_byte w 15 ->
    b16 = word_nth_byte w 16 ->
    b17 = word_nth_byte w 17 ->
    b18 = word_nth_byte w 18 ->
    b19 = word_nth_byte w 19 ->
    b20 = word_nth_byte w 20 ->
    b21 = word_nth_byte w 21 ->
    b22 = word_nth_byte w 22 ->
    b23 = word_nth_byte w 23 ->
    b24 = word_nth_byte w 24 ->
    b25 = word_nth_byte w 25 ->
    b26 = word_nth_byte w 26 ->
    b27 = word_nth_byte w 27 ->
    b28 = word_nth_byte w 28 ->
    b29 = word_nth_byte w 29 ->
    b30 = word_nth_byte w 30 ->
    b31 = word_nth_byte w 31 ->
    word_of_bytes
    [b0; b1; b2; b3; b4; b5; b6; b7; b8; b9; b10; b11; b12; b13; b14; b15; b16;
     b17; b18; b19; b20; b21; b22; b23; b24; b25; b26; b27; b28; b29; b30; b31] =
    w.
  Admitted.

  Axiom event : Set.

  Axiom memory_state : Set.
  Axiom empty_memory : memory_state.
  Axiom cut_memory : word -> word -> memory_state -> list byte.
  Axiom cut_memory_zero_nil :
    forall start m, cut_memory start word_zero m = nil.

  Module ST := FMapList.Make WordOrdered.

  Definition storage := ST.t word.

  Eval compute in ST.key.

  Definition storage_load (k : word) (m : storage) : word :=
    match ST.find k m with
    | None => word_zero
    | Some x => x
    end.
  Definition storage_store (k : WordOrdered.t) (v : word) (orig : storage) : storage :=
    if word_eq word_zero v then
      ST.remove k orig
    else
      ST.add k v orig.

  Definition empty_storage : storage := ST.empty word.
  Lemma empty_storage_empty : forall idx : WordOrdered.t,
      is_true (word_iszero (storage_load idx empty_storage)).
  Proof.
    intro idx.
    compute.
    auto.
  Qed.

  Lemma word_of_zero :
    word_zero = word_of_N 0.
  Proof.
    auto.
  Qed.
  Lemma word_of_one :
    word_one = word_of_N 1.
  Proof.
    auto.
  Qed.

  Definition word_of_nat :=
    BinInt.Z_of_nat.
End ConcreteWord.


Module ExamplesOnConcreteWord.

  Module ConcreteSem := (ContractSem.Make ConcreteWord).
  Include ConcreteSem.

  (** TODO: make this tactic only when immediate *)
  (** TODO: use this tactic *)
  Ltac compute_word_smaller :=
    set (focus := word_smaller _ _);
    compute in focus;
    unfold focus;
    clear focus.

  Ltac compute_word_mod :=
    set (focus := word_mod _ _);
    compute in focus;
    unfold focus;
    clear focus.

  Definition example2_program : program :=
    PUSH1 (word_of_N 0) ::
    SLOAD ::
    DUP1 ::
    PUSH1 (word_of_N 2) ::
    JUMPI ::
    PUSH1 (word_of_N 1) ::
    ADD ::
    PUSH1 (word_of_N 0) ::
    SSTORE ::
    PUSH1 (word_of_N 0) ::
    (* TODO: change some of these arguments to value, address *)
    PUSH1 (word_of_N 0) ::
    PUSH1 (word_of_N 0) ::
    PUSH1 (word_of_N 0) ::
    PUSH1 (word_of_N 0) ::
    PUSH1 (word_of_N 0) ::
    CALL ::
    ISZERO ::
    PUSH1 (word_of_N 0) ::
    JUMPI ::
    PUSH1 (word_of_N 0) ::
    PUSH1 (word_of_N 0) ::
    SSTORE ::
    STOP ::
    nil.

  Variable example2_address : address.

  Definition example2_depth_n_state  (n : word) (st : account_state) :=
    (n = 0%Z /\
       st.(account_address) = example2_address /\
       is_true (ST.equal word_eq (st.(account_storage)) empty_storage) /\
       st.(account_code) = example2_program /\
       st.(account_ongoing_calls) = nil ) \/
     (n = 1%Z /\
      st.(account_code) = example2_program /\
      storage_load 0%Z (account_storage st) = 1%Z /\
      st.(account_address) = example2_address /\
      is_true (ST.equal word_eq (storage_store 0%Z 0%Z st.(account_storage)) empty_storage)  /\
      exists ve, (st.(account_ongoing_calls) = ve :: nil /\
             ve.(venv_prg_sfx) =
    ISZERO ::
    PUSH1 (word_of_N 0) ::
    JUMPI ::
    PUSH1 (word_of_N 0) ::
    PUSH1 (word_of_N 0) ::
    SSTORE ::
    STOP ::
    nil
                  /\
                  is_true (ST.equal word_eq (storage_store 0%Z 0%Z ve.(venv_storage)) empty_storage) /\
   is_true (ST.equal word_eq (venv_storage_at_call ve) empty_storage))
     )
  .


Definition something_to_call :=
     {|
     callarg_gaslimit := 0%Z;
     callarg_code := address_of_word 0%Z;
     callarg_recipient := address_of_word 0%Z;
     callarg_value := 0%Z;
     callarg_data := cut_memory 0%Z 0%Z empty_memory;
     callarg_output_begin := 0%Z;
     callarg_output_size := storage_load 0%Z empty_storage |}.

(* TODO: remove duplicate somehow *)
CoFixpoint call_but_fail_on_reentrance (depth : word) :=
  if word_eq word_zero depth then
    Respond
      (fun _ =>
         ContractAction (ContractCall something_to_call)
              (call_but_fail_on_reentrance word_one))
      (fun _ => ContractAction ContractFail (call_but_fail_on_reentrance word_zero))
      (ContractAction ContractFail (call_but_fail_on_reentrance word_zero))
  else if word_eq word_one depth then
    Respond
      (fun _ => ContractAction ContractFail (call_but_fail_on_reentrance word_one))
      (fun _ => ContractAction (ContractReturn nil) (call_but_fail_on_reentrance word_zero))
      (ContractAction ContractFail (call_but_fail_on_reentrance word_zero))
  else
    Respond
      (fun _ => ContractAction ContractFail (call_but_fail_on_reentrance depth))
      (fun retval => ContractAction ContractFail (call_but_fail_on_reentrance (word_sub depth word_one)))
      (ContractAction ContractFail (call_but_fail_on_reentrance (word_sub depth word_one))).

  Lemma call_but_fail_on_reentrace_0_eq :
    call_but_fail_on_reentrance 0%Z =
    Respond
      (fun _ =>
         ContractAction (ContractCall something_to_call)
              (call_but_fail_on_reentrance word_one))
      (fun _ => ContractAction ContractFail (call_but_fail_on_reentrance word_zero))
      (ContractAction ContractFail (call_but_fail_on_reentrance word_zero)).
  Proof.
    rewrite (response_expander_eq (call_but_fail_on_reentrance 0%Z)).
    auto.
  Qed.

  Lemma call_but_fail_on_reentrace_1_eq :
    call_but_fail_on_reentrance 1%Z =
    Respond
      (fun _ => ContractAction ContractFail (call_but_fail_on_reentrance word_one))
      (fun retval => ContractAction (ContractReturn nil) (call_but_fail_on_reentrance word_zero))
      (ContractAction ContractFail (call_but_fail_on_reentrance word_zero)).
  Proof.
    rewrite (response_expander_eq (call_but_fail_on_reentrance 1%Z)).
    auto.
  Qed.

  Definition example2_spec (depth: word) : response_to_world :=
    call_but_fail_on_reentrance depth.

  Lemma update_remove_eq :
    forall orig,
      is_true (ST.equal word_eq orig empty_storage) ->
      is_true
        (ST.equal word_eq
                  (storage_store 0%Z 0%Z (ST.add 0%Z 1%Z orig))
                  empty_storage).
  Proof.
    intros orig nst2.
    apply ST.equal_1.
    split.
    {
      intro k.
      unfold storage_store.
      simpl.
      split.
      { intro H.
        apply False_ind.
        case_eq (word_eq k 0%Z).
        { intro k0.
          apply ST.Raw.remove_1 in H; auto.
          { apply ST.Raw.add_sorted.
            apply ST.sorted. }
          apply ST.E.eq_sym.
          assumption.
        }
        {
          intro neq.
          unfold ST.Raw.PX.In in H.
          case H as [e H].
          apply ST.Raw.remove_3 in H.
          {
            apply ST.Raw.add_3 in H.
            {
              apply ST.equal_2 in nst2.
              case nst2 as [I _].
              generalize (I k).
              unfold ST.Raw.PX.In.
              intro I'.
              case I' as [I0 _].
              simpl in I0.
              case I0.
              {
                exists e.
                apply H.
              }
              {
                intros x J.
                eapply ST.Raw.empty_1.
                apply J.
              }
            }
            {
              intro K.
              apply ST.E.eq_sym in K.
              congruence.
            }
          }
          {
            apply ST.Raw.add_sorted.
            apply ST.sorted.
          }
        }
      }
      {
        intro H.
        apply False_ind.
        case H.
        intros x Hx.
        apply (ST.Raw.empty_1 Hx).
      }
    }
    {
      intros k e e' H I.
      apply False_ind.
      generalize I.
      unfold empty_storage.
      generalize (ST.empty_1 I).
      auto.
    }
  Qed.

  Theorem example2_spec_impl_match :
    forall st n,
          example2_depth_n_state n st ->
          account_state_responds_to_world
            st (example2_spec n%Z) (fun _ _ => True).
  Proof.
    cofix.
    intros st n n_state.
    case n_state.
    {
      intro nst.
      destruct nst as [nst0 nst1].
      case nst1 as [nst1 nst2].
      case nst2 as [nst2 nst3].
      case nst3 as [nst3 nst4].
      subst.
      clear n_state.
      subst.
      unfold example2_spec.
      rewrite call_but_fail_on_reentrace_0_eq.
      apply AccountStep.
      {
        unfold respond_to_call_correctly.
        intros ce a con.
        split; [ solve [auto] | ].
        intros _ next.
        eexists.
        eexists.
        eexists.
        split.
        {
          intro s.
          simpl.
          rewrite nst3.
          repeat (case s as [| s]; [ solve [left; auto] | ]).
          assert (stl : forall idx, storage_load idx (account_storage st) = storage_load idx empty_storage).
          {
            intro idx.
            unfold storage_load.
            apply ST.equal_2 in nst2.
            unfold ST.Equivb in nst2.
            unfold ST.Raw.Equivb in nst2.
            simpl.
            case_eq (ST.find (elt:=word) idx (account_storage st)); auto.
            intros w H.
            apply ST.find_2 in H.
            apply False_ind.
            assert (ST.Raw.PX.In idx (ST.this (account_storage st))) as K.
            {
              unfold ST.Raw.PX.In.
              exists w.
              assumption.
            }
            case nst2 as [EE _].
            rewrite EE in K.
            unfold ST.Raw.PX.In in K.
            case K.
            intros content K'.
            apply (@ST.Raw.empty_1 word idx content).
            assumption.
          }
          simpl.
          rewrite !stl.
          unfold storage_load.
          unfold empty_storage.
          simpl.
          repeat (case s as [| s]; [ solve [left; auto] | ]).
          simpl.
          compute_word_mod.

          set (sm0 := word_smaller _ 0%Z).

          assert (H : sm0 = false).
          {
            unfold sm0.
            unfold word_smaller.
            simpl.
            rewrite ZModulo.spec_compare.
            set (v0 := (ZModulo.to_Z _ _)%Z).
            assert (0 <= v0)%Z.
            {
              apply (ZModulo.spec_to_Z_1).
              unfold ALEN.p.
              congruence.
            }
            set (comparison := (_ ?= _)%Z).
            case_eq comparison; try congruence.
            unfold comparison.
            rewrite Z.compare_nge_iff.
            intro H'.
            apply False_ind.
            apply H'.
            apply H.
          }
          rewrite H.

          right.
          f_equal.
          rewrite <- contract_action_expander_eq in next at 1.
          inversion next; subst.
          auto.
        }
        {
          simpl.
          rewrite <- contract_action_expander_eq in next at 1.
          inversion next; subst.
          simpl.
          apply example2_spec_impl_match.
          unfold example2_depth_n_state.
          right.
          split; auto.
          split; auto.
          split.
          {
            unfold storage_load.
            erewrite ST.find_1.
            { eauto. }
            apply ST.add_1.
            auto.
          }
          split; auto.
          split.
          {
            apply update_remove_eq.
            assumption.
          }
          eexists; eauto.
          split.
          {
            rewrite nst4.
            intuition.
          }
          {
            split; auto.
            split; auto.
            apply update_remove_eq.
            assumption.
          }

       (* this place should be come harder and harder as I specify the
           * state at depth 1
           *)
        }
      }
      {
        unfold respond_to_return_correctly.
        intros ? ? ? ?.
        simpl.
        rewrite nst4.
        congruence.
      }
      {
        intros ? ? ?.
        simpl.
        rewrite nst4.
        congruence.
      }
    }
    {
      intros H.
      destruct H as [n1 st_code].
      destruct st_code as [st_code st_load].
      destruct st_load as [st_load st_ongoing].
      subst.
      unfold example2_spec.
      rewrite call_but_fail_on_reentrace_1_eq.
      apply AccountStep.
      { (* call *)
        intros callenv act continuation.
        split; [solve [auto] | ].
        intros _ H.
        inversion H; subst.
        clear H.
        eexists.
        eexists.
        eexists.
        unfold build_venv_called.
        rewrite st_code.
        split.
        {
          intro s.
          repeat (case s as [| s]; [ solve [left; auto] | ]).

          simpl.
          compute_word_mod.
          unfold venv_first_instruction.
          rewrite st_load.
          simpl.
          rewrite st_code.
          simpl.
          right.
          eauto.
        }
        {
          apply example2_spec_impl_match.
          unfold example2_depth_n_state.
          intuition.
        }
      }
      { (* return *)
        unfold respond_to_return_correctly.
        intros rr venv cont act.
        elim st_ongoing.
        intros prev prevH.
        case prevH as [st_str prevH].
        case prevH as [prevH prevH'].
        case prevH' as [prevH' prevH''].
        case prevH'' as [prevH'' prevH'''].
        simpl.
        rewrite prevH'.
        intro H.
        inversion H; subst.
        clear H.
        intros act_cont_eq.
        eexists.
        eexists.
        eexists.
        split.
        {
          intro s.
          rewrite prevH''.
          repeat (case s as [| s]; [ solve [left; auto] | ]).
          simpl.
          right.
          f_equal.
          inversion act_cont_eq.
          auto.
        }
        {
          inversion act_cont_eq.
          apply example2_spec_impl_match.
          unfold example2_depth_n_state.
          left.
          repeat (split; auto); tauto.
        }
      }
      {
        unfold respond_to_fail_correctly.
        intros venv cont act.
        case st_ongoing as [st_addr st_ongoing].
        case st_ongoing as [st_storage st_ongoing].
        case st_ongoing as [ve veH].
        case veH as [st_ongoing ve_sfx].
        case ve_sfx as [ve_sfx ve_str].
        simpl.
        rewrite st_ongoing.
        intro venvH.
        inversion venvH; subst.
        clear venvH.
        intros act_cont_H.
        inversion act_cont_H; subst.
        clear act_cont_H.
        eexists.
        eexists.
        eexists.
        split.
        {
          intro s.
          rewrite ve_sfx.
          repeat (case s as [| s]; [ solve [left; auto] | ]).
          simpl.
          unfold compose.
          rewrite st_code.
          simpl.
          right.
          f_equal.
        }
        { (* update_account_state with contract_fail  *)
          simpl.
          apply example2_spec_impl_match.
          unfold example2_depth_n_state.
          left.
          repeat split; auto; tauto.
        }
      }
    }
  Qed.

  (** Example 4: a contract that keeps track of the accumulated income and spending.
   *
   * storage[0]: owner
   * storage[1]: income so far
   * storage[2]: spending so far
   * income so far - spending so far should coincide with the balance.
   *
   * data length 0 => receive eth; storage[1] should be incremented
   *
   * data length > 0 => not receiving eth
   * if msg.sender <> owner, abort.
   * data[0-19] is the address of recipient.
   * data[32-63] is the amount of spending.
   *
   * no particular prevention of re-entrancy.
   *)

  Definition failing_action cont : contract_behavior :=
    ContractAction ContractFail cont.

  Definition receive_eth cont : contract_behavior :=
    ContractAction (ContractReturn nil) cont.

  Definition sending_action (recipient : word) value cont : contract_behavior :=
    ContractAction (ContractCall
                      {|
                        callarg_gaslimit := 30000%Z;
                        callarg_code := address_of_word recipient;
                        callarg_recipient := address_of_word recipient;
                        callarg_value := value;
                        callarg_data := nil;
                        callarg_output_begin := 0%Z;
                        callarg_output_size := 0%Z
                      |}) cont.

  CoFixpoint counter_wallet (income_sofar : word) (spending_sofar : word)
    : response_to_world :=
    Respond
      (fun cenv =>
         match cenv.(callenv_data) with
         | nil => receive_eth (counter_wallet (word_add income_sofar cenv.(callenv_value)) spending_sofar)
         | _ =>
           if word_eq word_zero (cenv.(callenv_value)) then
             if Nat.leb 64 (List.length cenv.(callenv_data)) then
               let addr := list_slice 0 32 cenv.(callenv_data) in
               let value := list_slice 32 32 cenv.(callenv_data) in
               if word_smaller_or_eq value (word_sub (word_add income_sofar cenv.(callenv_value)) spending_sofar) then
                 sending_action addr value (counter_wallet income_sofar (word_add spending_sofar value))
               else
                 failing_action (counter_wallet income_sofar spending_sofar)
             else
               failing_action (counter_wallet income_sofar spending_sofar)
           else
             failing_action (counter_wallet income_sofar spending_sofar)
         end
      )
      (fun returned =>
         ContractAction (ContractReturn nil) (counter_wallet income_sofar spending_sofar)
      )
      (
        failing_action (counter_wallet income_sofar spending_sofar)
      ).

  Lemma counter_wallet_def :
    forall income_sofar spending_sofar,
      counter_wallet income_sofar spending_sofar =
    Respond
      (fun cenv =>
         match cenv.(callenv_data) with
         | nil => receive_eth (counter_wallet (word_add income_sofar cenv.(callenv_value)) spending_sofar)
         | _ =>
           if word_eq word_zero (cenv.(callenv_value)) then
             if Nat.leb 64 (List.length cenv.(callenv_data)) then
               let addr := list_slice 0 32 cenv.(callenv_data) in
               let value := list_slice 32 32 cenv.(callenv_data) in
               if word_smaller_or_eq value (word_sub (word_add income_sofar cenv.(callenv_value)) spending_sofar) then
                 sending_action addr value (counter_wallet income_sofar (word_add spending_sofar value))
               else
                 failing_action (counter_wallet income_sofar spending_sofar)
             else
               failing_action (counter_wallet income_sofar spending_sofar)
           else
             failing_action (counter_wallet income_sofar spending_sofar)
         end
      )
      (fun returned =>
         ContractAction (ContractReturn nil) (counter_wallet income_sofar spending_sofar)
      )
      (
        failing_action (counter_wallet income_sofar spending_sofar)
      ).
  Proof.
    intros i s.
    unfold counter_wallet.
    apply response_expander_eq.
  Qed.

  (* TODO: streamline this by allowing labels in JUMPDEST *)
  Definition plus_size_label : word := 13%Z.
  Arguments plus_size_label /.

  (* TODO: add owner as an immediate value and check it *)
  Definition counter_wallet_code : program :=
    CALLDATASIZE ::
      PUSH1 plus_size_label ::
        JUMPI ::
    (* size zero *)
    CALLVALUE ::
      PUSH1 word_zero (* storage[0] *) ::
        SLOAD ::
        ADD ::
      PUSH1 word_zero ::
        SSTORE ::
    STOP ::
    JUMPDEST (* plus_size_label *) ::
    CALLVALUE ::
      PUSH1 word_zero (* invalid destination *) ::
    (**) JUMPI ::
    (* call_value zero *)
    CALLDATASIZE ::
      PUSH1 (64%Z) ::
        instr_GT ::
      PUSH1 (0%Z) ::
        JUMPI (* data too small *) ::
    PUSH1 (0%Z) (* out size *) ::
      PUSH1 (0%Z) (* out offset *) ::
        PUSH1 (0%Z) (* out size *) ::
          PUSH1 (0%Z) (* in offset *) ::
            PUSH1 (0%Z) (* in size *) ::
              PUSH1 (32%Z) ::
                CALLDATALOAD (* value loaded *) ::
                DUP1 ::
                  PUSH1 (1%Z) ::
                    SLOAD ::
                    ADD ::
                  PUSH1 (1%Z) ::
                    SSTORE ::
                PUSH1 (0%Z) ::
                  CALLDATALOAD (* addr loaded *) ::
                  PUSH2 (30000%Z) ::
                    CALL ::
      ISZERO ::
      PUSH1 word_zero ::
        JUMPI ::
    STOP ::
    nil.


  Definition counter_wallet_invariant (v : variable_env) (c : constant_env) : Prop :=
      word_add (v.(venv_balance) c.(cenv_this)) (storage_load 1%Z v.(venv_storage))
    = word_add v.(venv_value_sent) (storage_load 0%Z v.(venv_storage)).

  Axiom counter_wallet_address : address.

  Definition counter_wallet_storage (income_sofar spending_sofar : word) : storage :=
    storage_store 1%Z spending_sofar (storage_store 0%Z income_sofar (ST.empty word))
    .

  Definition counter_wallet_account_state (income_sofar spending_sofar : word) (going_calls : list variable_env) : account_state :=
    {|
      account_address := counter_wallet_address (* TODO: declare this in a section *);
      account_storage := counter_wallet_storage income_sofar spending_sofar ;
      account_code := counter_wallet_code ;
      account_balance := word_sub income_sofar spending_sofar ;
      account_ongoing_calls := going_calls
    |}
    .

  Record counter_wallet_calling_state (v : variable_env) :=
    {
      cw_calling_prg_sfx :
        (v.(venv_prg_sfx) =
         ISZERO ::
             PUSH1 word_zero ::
             JUMPI ::
             STOP ::
             nil)
    }.

  Definition all_cw_calling_state lst :=
    forall v, In v lst -> counter_wallet_calling_state v.

  Lemma all_cw_calling_state_head_tail :
    forall head tail,
      all_cw_calling_state (head :: tail) ->
      all_cw_calling_state tail /\ counter_wallet_calling_state head.
  Proof.
    intros head tail H.
    split.
    {
      intro elm.
      intro elmh.
      apply H.
      apply in_cons.
      auto.
    }
    apply H.
    apply in_eq.
  Qed.

  Theorem counter_wallet_correct :
    forall (income_sofar spending_sofar : word) ongoing,
      all_cw_calling_state ongoing ->
      account_state_responds_to_world
        (counter_wallet_account_state income_sofar spending_sofar ongoing)
        (counter_wallet income_sofar spending_sofar)
        counter_wallet_invariant.
    (* TODO: strengthen the statement so that coinduction goes through. *)
  Proof.
    cofix.
    intros income_sofar spending_sofar ongoing ongoingH.
    rewrite counter_wallet_def.
    apply AccountStep.
    {
      unfold respond_to_call_correctly.
      intros callenv act cont.
      split.
      {
        unfold counter_wallet_invariant.
        simpl.
        unfold update_balance.
        rewrite address_eq_refl.
        unfold counter_wallet_storage.
        set (spend := storage_load 1%Z _).
        (* TODO: a geneeral lemma is needed here *)
        assert (spendH : spend = spending_sofar) by admit.
        rewrite spendH.
        set (income := storage_load 0%Z _).
        assert (incomeH : income = income_sofar) by admit.
        rewrite incomeH.
        rewrite !addsub.
        rewrite addK.
        apply addC.
      }
      {
        intro I.
        case_eq (callenv_data callenv).
        { (* input data is nil *)
          intro data_nil.
          unfold receive_eth.
          intro H.
          inversion H; subst.
          clear H.
          eexists.
          eexists.
          eexists.
          split.
          {
            intro s.
            repeat (case s as [| s]; [ solve [left; auto] | cbn ]).
            rewrite data_nil.
            repeat (case s as [| s]; [ solve [left; auto] | cbn ]).
            right.
            reflexivity.
          }
          {
            cbn.
            unfold counter_wallet_storage.
            unfold storage_load.
            unfold ZModulo.zero.
            set (prev_income := ST.find _ _).
            assert (P : prev_income = Some income_sofar) by admit.
            rewrite P.
            set (new_income := ZModulo.add income_sofar _).
            generalize (counter_wallet_correct new_income).
            intro IH.
            unfold counter_wallet_account_state in IH.
            unfold counter_wallet_storage in IH.
            assert (II : storage_store 0%Z new_income
                         (storage_store 1%Z spending_sofar
                            (storage_store 0%Z income_sofar
                               (ST.empty word))) =
                         (storage_store 1%Z spending_sofar
                            (storage_store 0%Z new_income
                               (ST.empty word)))) by admit.
            rewrite II.
            unfold update_balance.
            rewrite address_eq_refl.
            rewrite addsub.
            eapply IH.
            assumption.
          }
        }
        { (* input data is not nil *)
          intros b l bl_eq.
          case_eq (word_eq word_zero (callenv_value callenv)).
          { (* sent value is zero *)
            intro sent_zero.
            (* hmmm wanting ssreflect tactics. *)
            match goal with
              | [ |- ((if ?t then _ else _) = _) -> _] => case_eq t
            end.
            {
              intro data_big_enough.
              unfold sending_action.
              (* Here, before introducing the existential variables,
               * all ambuiguities must be resolved. *)
              set (enough_balance_spec := word_smaller_or_eq _ _).
              case_eq enough_balance_spec.
              { (* enough balance *)
                intro enough_balance_spec_t.
                intro H.
                inversion H; subst.
                clear H.
                eexists.
                eexists.
                eexists.
                split.
                {
                  intro s.
                  repeat (case s as [| s]; [ solve [left; auto] | ]).
                  cbn.
                  unfold datasize.
                  cbn.
                  set (e0 := ZModulo.eq0 _ _).
                  assert (R : e0 = false) by admit.
                  rewrite R.
                  unfold N_of_word.
                  cbn.
                  unfold ZModulo.to_Z.
                  unfold ZModulo.wB.
                  simpl.
                  repeat (case s as [| s]; [ solve [left; auto] | ]).
                  simpl.
                  assert (Z : word_iszero (callenv_value callenv) = true) by admit.
                  rewrite Z.
                  repeat (case s as [| s]; [ solve [left; auto] | ]).
                  cbn.
                  unfold datasize.
                  cbn.
                  set (s64 := word_smaller _ _).
                  assert (S : s64 = false) by admit.
                  rewrite S.
                  simpl.
                  repeat (case s as [| s]; [ solve [left; auto] | cbn ]).
                  set (balance_smaller := word_smaller _ _).
                  assert (F : balance_smaller = false)by admit (* use enough_balance_spec *).
                  rewrite F.
                  clear F.
                  right.
                  f_equal.
                  f_equal.
                  f_equal.
                  {
                    unfold cut_data.
                    simpl.
                    rewrite bl_eq.
                    reflexivity.
                  }
                  {
                    unfold cut_data.
                    simpl.
                    rewrite bl_eq.
                    reflexivity.
                  }
                  {
                    unfold cut_data.
                    simpl.
                    rewrite bl_eq.
                    reflexivity.
                  }
                  {
                    (* TODO: need to define cut_memory *)
                    admit.
                  }
                }
                {
                  cbn.
                  unfold cut_data.
                  cbn.
                  unfold counter_wallet_account_state in counter_wallet_correct.
                  set (new_storage := storage_store _ _ _).
                  set (new_ongoing := _ :: ongoing).
                  unfold update_balance.
                  rewrite address_eq_refl.
                  set (new_balance := if (_ : bool) then _ else _).
                  set (new_sp := ZModulo.add spending_sofar _).
                  assert (S : new_storage = counter_wallet_storage income_sofar new_sp) by admit.
                  rewrite S.
                  assert (B : new_balance = word_sub income_sofar new_sp) by admit.
                  rewrite B.
                  apply (counter_wallet_correct income_sofar new_sp).
                  unfold new_ongoing.
                  unfold all_cw_calling_state.
                  intros elm elmH.
                  apply in_inv in elmH.
                  case elmH.
                  {
                    intro K.
                    rewrite <-K.
                    apply Build_counter_wallet_calling_state.
                    reflexivity.
                  }
                  {
                    apply ongoingH.
                  }
                }
              }
              { (* not enough balance *)
                intro not_enough_spec.
                intro H.
                inversion H; subst.
                clear H.

                eexists.
                eexists.
                eexists.
                split.
                {
                  intro s.
                  repeat (case s as [| s]; [ solve [left; auto] | ]).
                  cbn.
                  unfold datasize.
                  cbn.
                  set (e0 := ZModulo.eq0 _ _).
                  assert (R : e0 = false) by admit.
                  rewrite R.
                  unfold N_of_word.
                  cbn.
                  unfold ZModulo.to_Z.
                  unfold ZModulo.wB.
                  simpl.
                  repeat (case s as [| s]; [ solve [left; auto] | ]).
                  simpl.
                  assert (Z : word_iszero (callenv_value callenv) = true) by admit.
                  rewrite Z.
                  repeat (case s as [| s]; [ solve [left; auto] | ]).
                  cbn.
                  unfold datasize.
                  simpl.
                  set (s64 := word_smaller _ _).
                  assert (S : s64 = false) by admit.
                  rewrite S.
                  simpl.
                  repeat (case s as [| s]; [ solve [left; auto] | cbn ]).
                  set (cd := cut_data _ _).
                  assert (cdH : cd = list_slice 0 32 (callenv_data callenv)) by admit.
                  rewrite cdH.
                  clear cdH cd.
                  set (balance_smaller := word_smaller _ _).
                  assert (A : balance_smaller = true) by admit.
                  rewrite A.
                  right.
                  eauto.
                }
                {
                  simpl.
                  unfold counter_wallet_account_state in counter_wallet_correct.
                  unfold update_balance.
                  rewrite address_eq_refl.
                  apply counter_wallet_correct.
                  assumption.
                }
              }
            }
            {
              intro data_short.
              unfold failing_action.
              intro H.
              inversion H; subst.
              clear H.
              eexists.
              eexists.
              eexists.
              split.
              {
                intros s.
                repeat (case s as [| s]; [ solve [left; auto] | cbn ]).
                unfold plus_size_label.
                unfold datasize.
                cbn.
                set (zero_cond := ZModulo.eq0 _ _ ).
                assert (Zf : zero_cond = false) by admit.
                rewrite Zf.
                cbn.
                simpl.
                repeat (case s as [| s]; [ solve [left; auto] | ]).
                cbn.
                set (z_cond := ZModulo.eq0 _ _).
                assert (Zt : z_cond = true) by admit.
                rewrite Zt.
                repeat (case s as [| s]; [ solve [left; auto] | ]).
                cbn.
                unfold datasize.
                cbn.
                set (small := word_smaller _ _).
                assert (SS : small = true) by admit.
                rewrite SS.
                simpl.
                right.
                eauto.
              }
              {
                unfold update_account_state.
                cbn.
                unfold update_balance.
                rewrite address_eq_refl.
                apply counter_wallet_correct.
                assumption.
              }
            }
          }
          { (* sent value is not zero, and data is also sent; should fail *)
            (* I can just imagine this needs the definition of datasize, too *)
            idtac.
            intro value_nonzero.
            intro H.
            inversion H; subst.
            eexists.
            eexists.
            eexists.
            split.
            {
              intro s.
              repeat (case s as [| s]; [ solve [left; auto] | ]).
              cbn.
              unfold datasize.
              cbn.
              set (e0 := ZModulo.eq0 _ _).
              assert (E0 : e0 = false) by admit (* an extra assumption that data is not as long as 2^256 is needed*).
              rewrite E0.
              simpl.
              (* TODO: define a lemma so that just proving something for a large s is enough *)
              repeat (case s as [| s]; [ solve [left; auto] | ]).
              cbn.
              set (v0 := ZModulo.eq0 _ _).
              assert (V0 : v0 = false) by admit.
              rewrite V0.
              cbn.
              right. (* TODO: maybe name a constructor *)
              eauto.
            }
            {
                unfold update_account_state.
                cbn.
                unfold update_balance.
                rewrite address_eq_refl.
                apply counter_wallet_correct.
                assumption.
            }
          }
        }
      }
    }
    {
      (* Now this goal does make sense *)
      (* TODO: maybe try to see the required condition here? *)
      unfold respond_to_return_correctly.
      intros rr venv cont act.
      intro venvH.
      intro H.
      inversion H; subst.
      clear H.
      unfold build_venv_returned in venvH.
      unfold counter_wallet_account_state in venvH.
      cbn in venvH.
      case ongoing as [| recovered rest_oging]; try congruence.
      (* TODO: define a property that implies this goal *)
      eexists.
      eexists.
      eexists.
      split.
      {
        inversion venvH; subst.
        clear venvH.
        unfold all_cw_calling_state in ongoingH.
        assert (CSR : counter_wallet_calling_state recovered)
          by (* TODO: use all_cw_calling_state *) admit.
        rewrite (cw_calling_prg_sfx _ CSR).
        intro s.
        repeat (case s as [| s]; [ solve [left; auto] | ]).
        simpl.
        right.
        f_equal.
        }
      {
        unfold update_account_state.
        unfold counter_wallet_account_state in counter_wallet_correct.
        unfold account_state_update_storage.
        simpl.

        rewrite get_update_balance.
        apply counter_wallet_correct.


        apply all_cw_calling_state_head_tail in ongoingH.
        tauto.
      }
    }
    {
      unfold respond_to_fail_correctly.
      intros v c a.
      intro v_eq.
      intro a_c_eq.
      inversion a_c_eq; subst.
      unfold failing_action in a_c_eq.
      clear a_c_eq.
      unfold build_venv_fail in v_eq.
      simpl in v_eq.
      case_eq ongoing.
      {
        intros ?.
        subst.
        congruence.
      }
      intros ongoing_head ongoing_tail ongoing_eq.
      subst.
      inversion v_eq; subst.
      clear v_eq.
      eexists.
      eexists.
      eexists.
      split.
      {
        intro s.
        repeat (case s as [| s]; [ solve [left; auto] | cbn ]).

        admit.
      }
      {
        admit.
      }
    }
  Admitted.

End ExamplesOnConcreteWord.

(* TODO: currently,
   lack of balance is treated in the semantics, but lack of gas is not.
   This discrepancy needs to be solved.
*)
